--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:49:27 05/19/2021
-- Design Name:   
-- Module Name:   /mnt/e/JU/8/VLSI/Lab/Code/Assignment7/TFlipflopDownCounterTestBench.vhd
-- Project Name:  Assignment7
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: TFlipflopDownCounter
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY TFlipflopDownCounterTestBench IS
END TFlipflopDownCounterTestBench;
 
ARCHITECTURE behavior OF TFlipflopDownCounterTestBench IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT TFlipflopDownCounter
    PORT(
         rst : IN  std_logic;
         clk : IN  std_logic;
         qqqq : INOUT  std_logic_vector(2 downto 0);
         qqqqbar : INOUT  std_logic_vector(2 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal rst : std_logic := '0';
   signal clk : std_logic := '0';

	--BiDirs
   signal qqqq : std_logic_vector(2 downto 0);
   signal qqqqbar : std_logic_vector(2 downto 0);

   -- Clock period definitions
   --constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: TFlipflopDownCounter PORT MAP (
          rst => rst,
          clk => clk,
          qqqq => qqqq,
          qqqqbar => qqqqbar
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for 1 ps;
		clk <= '1';
		wait for 1 ps;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      rst<='0';
		wait for 1 ps;
		rst<='1';
		wait for 1 ps;
		rst<='0';
		wait for 1 ps;
		loop1:loop
			wait for 1 ps;
			wait for 1 ps;
		end loop;
   end process;

END;
